magic
tech scmos
timestamp 1543430412
<< polysilicon >>
rect 14 213 18 219
rect 196 214 200 220
rect 14 187 18 193
rect 96 187 100 203
rect 196 188 200 194
rect 278 188 282 204
rect 14 171 18 177
rect 14 111 18 161
rect 96 111 100 177
rect 196 172 200 178
rect 14 107 28 111
rect 40 107 44 111
rect 62 107 66 111
rect 86 107 100 111
rect 14 35 18 107
rect 96 35 100 107
rect 14 31 28 35
rect 48 31 52 35
rect 68 31 72 35
rect 84 31 100 35
rect 196 112 200 162
rect 278 112 282 178
rect 196 108 210 112
rect 222 108 226 112
rect 244 108 248 112
rect 268 108 282 112
rect 196 36 200 108
rect 278 36 282 108
rect 196 32 210 36
rect 230 32 234 36
rect 250 32 254 36
rect 266 32 282 36
rect 14 -36 18 31
rect 96 -36 100 31
rect 14 -40 28 -36
rect 40 -40 45 -36
rect 60 -40 66 -36
rect 86 -40 100 -36
rect 14 -122 18 -40
rect 96 -122 100 -40
rect 14 -126 28 -122
rect 48 -126 52 -122
rect 70 -126 74 -122
rect 86 -126 100 -122
<< ndiffusion >>
rect -8 161 -6 171
rect 4 161 14 171
rect 18 161 28 171
rect 38 161 40 171
rect 28 131 40 133
rect 28 111 40 119
rect 174 162 176 172
rect 186 162 196 172
rect 200 162 210 172
rect 220 162 222 172
rect 28 99 40 107
rect 28 85 40 87
rect 72 55 84 57
rect 72 35 84 43
rect 210 132 222 134
rect 210 112 222 120
rect 210 100 222 108
rect 210 86 222 88
rect 254 56 266 58
rect 254 36 266 44
rect 72 23 84 31
rect 72 9 84 11
rect 28 -15 40 -13
rect 28 -36 40 -27
rect 254 24 266 32
rect 254 10 266 12
rect 28 -47 40 -40
rect 28 -61 40 -59
rect 74 -101 86 -99
rect 74 -122 86 -113
rect 74 -133 86 -126
rect 74 -147 86 -145
<< pdiffusion >>
rect -8 209 14 213
rect -8 199 -6 209
rect 4 199 14 209
rect -8 193 14 199
rect 18 209 40 213
rect 18 199 28 209
rect 38 199 40 209
rect 174 210 196 214
rect 18 193 40 199
rect 174 200 176 210
rect 186 200 196 210
rect 174 194 196 200
rect 200 210 222 214
rect 200 200 210 210
rect 220 200 222 210
rect 200 194 222 200
rect 66 131 86 133
rect 66 119 70 131
rect 82 119 86 131
rect 66 111 86 119
rect 66 99 86 107
rect 66 87 70 99
rect 82 87 86 99
rect 66 85 86 87
rect 28 55 48 57
rect 28 43 32 55
rect 44 43 48 55
rect 28 35 48 43
rect 248 132 268 134
rect 248 120 252 132
rect 264 120 268 132
rect 248 112 268 120
rect 248 100 268 108
rect 248 88 252 100
rect 264 88 268 100
rect 248 86 268 88
rect 210 56 230 58
rect 210 44 214 56
rect 226 44 230 56
rect 210 36 230 44
rect 28 23 48 31
rect 28 11 32 23
rect 44 11 48 23
rect 28 9 48 11
rect 66 -15 86 -13
rect 66 -27 70 -15
rect 82 -27 86 -15
rect 66 -36 86 -27
rect 210 24 230 32
rect 210 12 214 24
rect 226 12 230 24
rect 210 10 230 12
rect 66 -47 86 -40
rect 66 -59 70 -47
rect 82 -59 86 -47
rect 66 -61 86 -59
rect 28 -101 48 -99
rect 28 -113 32 -101
rect 44 -113 48 -101
rect 28 -122 48 -113
rect 28 -133 48 -126
rect 28 -145 32 -133
rect 44 -145 48 -133
rect 28 -147 48 -145
<< metal1 >>
rect -6 224 186 233
rect -6 209 4 224
rect 176 210 186 224
rect 28 187 38 199
rect 210 188 220 200
rect 2 177 8 187
rect 28 177 90 187
rect 184 178 190 188
rect 210 178 272 188
rect 28 171 38 177
rect 210 172 220 178
rect -6 153 4 161
rect 176 153 186 162
rect -6 145 186 153
rect -10 119 28 131
rect 40 119 70 131
rect 162 120 210 132
rect 222 120 252 132
rect 40 87 70 99
rect 52 75 62 87
rect 162 75 172 120
rect 222 88 252 100
rect 52 65 172 75
rect 234 76 244 88
rect 234 66 294 76
rect 52 55 62 65
rect 234 56 244 66
rect 44 43 72 55
rect 226 44 254 56
rect -10 11 32 23
rect 44 11 72 23
rect 166 12 214 24
rect 226 12 254 24
rect -10 -26 28 -15
rect 40 -27 70 -15
rect 40 -59 70 -47
rect 52 -76 61 -59
rect 166 -76 178 12
rect 52 -84 178 -76
rect 52 -101 61 -84
rect 44 -113 74 -101
rect -13 -145 32 -133
rect 44 -145 74 -133
<< ntransistor >>
rect 14 161 18 171
rect 196 162 200 172
rect 28 107 40 111
rect 72 31 84 35
rect 210 108 222 112
rect 254 32 266 36
rect 28 -40 40 -36
rect 74 -126 86 -122
<< ptransistor >>
rect 14 193 18 213
rect 196 194 200 214
rect 66 107 86 111
rect 28 31 48 35
rect 248 108 268 112
rect 210 32 230 36
rect 66 -40 86 -36
rect 28 -126 48 -122
<< polycontact >>
rect 8 177 18 187
rect 90 177 100 187
rect 190 178 200 188
rect 272 178 282 188
<< ndcontact >>
rect -6 161 4 171
rect 28 161 38 171
rect 28 119 40 131
rect 176 162 186 172
rect 210 162 220 172
rect 28 87 40 99
rect 72 43 84 55
rect 210 120 222 132
rect 210 88 222 100
rect 254 44 266 56
rect 72 11 84 23
rect 28 -27 40 -15
rect 254 12 266 24
rect 28 -59 40 -47
rect 74 -113 86 -101
rect 74 -145 86 -133
<< pdcontact >>
rect -6 199 4 209
rect 28 199 38 209
rect 176 200 186 210
rect 210 200 220 210
rect 70 119 82 131
rect 70 87 82 99
rect 32 43 44 55
rect 252 120 264 132
rect 252 88 264 100
rect 214 44 226 56
rect 32 11 44 23
rect 70 -27 82 -15
rect 214 12 226 24
rect 70 -59 82 -47
rect 32 -113 44 -101
rect 32 -145 44 -133
<< labels >>
rlabel metal1 -2 219 -2 219 5 Vdd
rlabel metal1 -2 147 -2 147 1 GND
rlabel metal1 -6 125 -6 125 3 Input1
rlabel metal1 -6 17 -6 17 3 Input2
rlabel metal1 180 220 180 220 5 Vdd
rlabel metal1 180 148 180 148 1 GND
rlabel metal1 290 70 290 70 7 Output
rlabel metal1 5 182 5 182 1 Ctrl1
rlabel metal1 186 183 186 183 1 Ctrl2
rlabel metal1 -4 -21 -4 -21 1 Input3
rlabel metal1 -7 -139 -7 -139 1 Input4
<< end >>

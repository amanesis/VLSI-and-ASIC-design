magic
tech scmos
timestamp 1543609882
<< polysilicon >>
rect 122 1013 126 1020
rect 12 970 19 979
rect 54 960 58 980
rect 122 960 126 1008
rect 412 988 416 994
rect 194 956 198 976
rect 412 962 416 968
rect 494 962 498 978
rect 54 916 58 940
rect 122 916 126 940
rect 412 946 416 952
rect 194 930 198 936
rect 270 930 274 942
rect 194 914 198 920
rect 54 860 58 906
rect 122 860 126 906
rect 194 898 198 904
rect 202 858 206 878
rect 270 858 274 920
rect 412 886 416 936
rect 494 886 498 952
rect 412 882 426 886
rect 438 882 442 886
rect 460 882 464 886
rect 484 882 498 886
rect 54 816 58 840
rect 122 816 126 840
rect 202 834 206 838
rect 202 814 206 824
rect 270 814 274 838
rect 302 831 306 837
rect 54 786 58 806
rect 122 786 126 806
rect 202 784 206 804
rect 270 784 274 804
rect 302 749 306 824
rect 412 810 416 882
rect 494 810 498 882
rect 547 850 551 863
rect 412 806 426 810
rect 446 806 450 810
rect 466 806 470 810
rect 482 806 498 810
rect 394 777 402 790
rect 135 687 139 749
rect 203 745 306 749
rect 203 687 207 745
rect 479 689 483 709
rect 547 689 551 840
rect 815 731 819 733
rect 325 679 329 685
rect 135 643 139 667
rect 203 643 207 667
rect 669 681 673 687
rect 325 653 329 659
rect 479 645 483 669
rect 547 645 551 669
rect 669 655 673 661
rect 325 637 329 643
rect 88 600 96 606
rect 135 533 139 633
rect 203 533 207 633
rect 669 639 673 645
rect 325 621 329 627
rect 275 529 279 549
rect 479 535 483 635
rect 547 535 551 635
rect 669 623 673 629
rect 815 613 819 721
rect 1033 659 1037 685
rect 883 613 887 633
rect 993 617 997 623
rect 815 569 819 593
rect 883 569 887 593
rect 993 591 997 597
rect 993 575 997 581
rect 993 559 997 565
rect 135 489 139 513
rect 203 489 207 513
rect 619 531 623 551
rect 815 539 819 559
rect 883 537 887 559
rect 275 503 279 509
rect 351 503 355 515
rect 275 487 279 493
rect 135 433 139 479
rect 203 433 207 479
rect 275 471 279 477
rect 283 431 287 451
rect 351 431 355 493
rect 479 491 483 515
rect 547 491 551 515
rect 883 525 887 527
rect 619 505 623 511
rect 695 505 699 517
rect 619 489 623 495
rect 479 435 483 481
rect 547 435 551 481
rect 619 473 623 479
rect 135 389 139 413
rect 203 389 207 413
rect 627 433 631 453
rect 695 433 699 495
rect 283 407 287 411
rect 283 387 287 397
rect 351 387 355 411
rect 479 403 483 415
rect 389 399 483 403
rect 479 391 483 399
rect 547 391 551 415
rect 627 409 631 413
rect 135 359 139 379
rect 203 359 207 379
rect 627 389 631 399
rect 695 389 699 413
rect 733 401 747 405
rect 283 357 287 377
rect 351 357 355 377
rect 479 361 483 381
rect 547 361 551 381
rect 627 359 631 379
rect 695 359 699 379
<< ndiffusion >>
rect 390 936 392 946
rect 402 936 412 946
rect 416 936 426 946
rect 436 936 438 946
rect 36 906 38 916
rect 48 906 54 916
rect 58 906 122 916
rect 126 906 130 916
rect 140 906 142 916
rect 172 904 174 914
rect 184 904 194 914
rect 198 904 208 914
rect 218 904 220 914
rect 426 906 438 908
rect 426 886 438 894
rect 36 806 38 816
rect 48 806 54 816
rect 58 806 80 816
rect 90 806 122 816
rect 126 806 130 816
rect 140 806 142 816
rect 184 804 186 814
rect 196 804 202 814
rect 206 804 228 814
rect 238 804 270 814
rect 274 804 278 814
rect 288 804 290 814
rect 426 874 438 882
rect 426 860 438 862
rect 470 830 482 832
rect 470 810 482 818
rect 470 798 482 806
rect 470 784 482 786
rect 117 633 119 643
rect 129 633 135 643
rect 139 633 203 643
rect 207 633 211 643
rect 221 633 223 643
rect 303 627 305 637
rect 315 627 325 637
rect 329 627 339 637
rect 349 627 351 637
rect 461 635 463 645
rect 473 635 479 645
rect 483 635 547 645
rect 551 635 555 645
rect 565 635 567 645
rect 647 629 649 639
rect 659 629 669 639
rect 673 629 683 639
rect 693 629 695 639
rect 797 559 799 569
rect 809 559 815 569
rect 819 559 841 569
rect 851 559 883 569
rect 887 559 891 569
rect 901 559 903 569
rect 971 565 973 575
rect 983 565 993 575
rect 997 565 1007 575
rect 1017 565 1019 575
rect 117 479 119 489
rect 129 479 135 489
rect 139 479 203 489
rect 207 479 211 489
rect 221 479 223 489
rect 253 477 255 487
rect 265 477 275 487
rect 279 477 289 487
rect 299 477 301 487
rect 461 481 463 491
rect 473 481 479 491
rect 483 481 547 491
rect 551 481 555 491
rect 565 481 567 491
rect 597 479 599 489
rect 609 479 619 489
rect 623 479 633 489
rect 643 479 645 489
rect 117 379 119 389
rect 129 379 135 389
rect 139 379 161 389
rect 171 379 203 389
rect 207 379 211 389
rect 221 379 223 389
rect 265 377 267 387
rect 277 377 283 387
rect 287 377 309 387
rect 319 377 351 387
rect 355 377 359 387
rect 369 377 371 387
rect 461 381 463 391
rect 473 381 479 391
rect 483 381 505 391
rect 515 381 547 391
rect 551 381 555 391
rect 565 381 567 391
rect 609 379 611 389
rect 621 379 627 389
rect 631 379 653 389
rect 663 379 695 389
rect 699 379 703 389
rect 713 379 715 389
<< pdiffusion >>
rect 390 984 412 988
rect 36 954 54 960
rect 36 944 38 954
rect 48 944 54 954
rect 36 940 54 944
rect 58 954 122 960
rect 58 944 80 954
rect 90 944 122 954
rect 58 940 122 944
rect 126 954 142 960
rect 390 974 392 984
rect 402 974 412 984
rect 390 968 412 974
rect 416 984 438 988
rect 416 974 426 984
rect 436 974 438 984
rect 416 968 438 974
rect 126 944 130 954
rect 140 944 142 954
rect 126 940 142 944
rect 172 952 194 956
rect 172 942 174 952
rect 184 942 194 952
rect 172 936 194 942
rect 198 952 220 956
rect 198 942 208 952
rect 218 942 220 952
rect 198 936 220 942
rect 36 854 54 860
rect 36 844 38 854
rect 48 844 54 854
rect 36 840 54 844
rect 58 840 122 860
rect 126 854 142 860
rect 464 906 484 908
rect 464 894 468 906
rect 480 894 484 906
rect 464 886 484 894
rect 126 844 130 854
rect 140 844 142 854
rect 126 840 142 844
rect 184 852 202 858
rect 184 842 186 852
rect 196 842 202 852
rect 184 838 202 842
rect 206 838 270 858
rect 274 852 290 858
rect 274 842 278 852
rect 288 842 290 852
rect 274 838 290 842
rect 464 874 484 882
rect 464 862 468 874
rect 480 862 484 874
rect 464 860 484 862
rect 426 830 446 832
rect 426 818 430 830
rect 442 818 446 830
rect 426 810 446 818
rect 426 798 446 806
rect 426 786 430 798
rect 442 786 446 798
rect 426 784 446 786
rect 117 681 135 687
rect 117 671 119 681
rect 129 671 135 681
rect 117 667 135 671
rect 139 681 203 687
rect 139 671 161 681
rect 171 671 203 681
rect 139 667 203 671
rect 207 681 223 687
rect 207 671 211 681
rect 221 671 223 681
rect 461 683 479 689
rect 207 667 223 671
rect 303 675 325 679
rect 303 665 305 675
rect 315 665 325 675
rect 303 659 325 665
rect 329 675 351 679
rect 329 665 339 675
rect 349 665 351 675
rect 461 673 463 683
rect 473 673 479 683
rect 461 669 479 673
rect 483 683 547 689
rect 483 673 505 683
rect 515 673 547 683
rect 483 669 547 673
rect 551 683 567 689
rect 551 673 555 683
rect 565 673 567 683
rect 551 669 567 673
rect 647 677 669 681
rect 329 659 351 665
rect 647 667 649 677
rect 659 667 669 677
rect 647 661 669 667
rect 673 677 695 681
rect 673 667 683 677
rect 693 667 695 677
rect 673 661 695 667
rect 117 527 135 533
rect 117 517 119 527
rect 129 517 135 527
rect 117 513 135 517
rect 139 527 203 533
rect 139 517 161 527
rect 171 517 203 527
rect 139 513 203 517
rect 207 527 223 533
rect 971 613 993 617
rect 797 607 815 613
rect 797 597 799 607
rect 809 597 815 607
rect 797 593 815 597
rect 819 593 883 613
rect 887 607 903 613
rect 887 597 891 607
rect 901 597 903 607
rect 971 603 973 613
rect 983 603 993 613
rect 971 597 993 603
rect 997 613 1019 617
rect 997 603 1007 613
rect 1017 603 1019 613
rect 997 597 1019 603
rect 887 593 903 597
rect 461 529 479 535
rect 207 517 211 527
rect 221 517 223 527
rect 207 513 223 517
rect 253 525 275 529
rect 253 515 255 525
rect 265 515 275 525
rect 253 509 275 515
rect 279 525 301 529
rect 279 515 289 525
rect 299 515 301 525
rect 461 519 463 529
rect 473 519 479 529
rect 461 515 479 519
rect 483 529 547 535
rect 483 519 505 529
rect 515 519 547 529
rect 483 515 547 519
rect 551 529 567 535
rect 551 519 555 529
rect 565 519 567 529
rect 551 515 567 519
rect 597 527 619 531
rect 597 517 599 527
rect 609 517 619 527
rect 279 509 301 515
rect 117 427 135 433
rect 117 417 119 427
rect 129 417 135 427
rect 117 413 135 417
rect 139 413 203 433
rect 207 427 223 433
rect 597 511 619 517
rect 623 527 645 531
rect 623 517 633 527
rect 643 517 645 527
rect 623 511 645 517
rect 207 417 211 427
rect 221 417 223 427
rect 207 413 223 417
rect 265 425 283 431
rect 265 415 267 425
rect 277 415 283 425
rect 265 411 283 415
rect 287 411 351 431
rect 355 425 371 431
rect 355 415 359 425
rect 369 415 371 425
rect 461 429 479 435
rect 461 419 463 429
rect 473 419 479 429
rect 461 415 479 419
rect 483 415 547 435
rect 551 429 567 435
rect 551 419 555 429
rect 565 419 567 429
rect 551 415 567 419
rect 609 427 627 433
rect 609 417 611 427
rect 621 417 627 427
rect 355 411 371 415
rect 609 413 627 417
rect 631 413 695 433
rect 699 427 715 433
rect 699 417 703 427
rect 713 417 715 427
rect 699 413 715 417
<< metal1 >>
rect 127 1008 146 1013
rect 300 993 402 1001
rect 300 972 310 993
rect 392 984 402 993
rect 2 970 310 972
rect 2 965 12 970
rect 19 965 310 970
rect 2 962 310 965
rect 426 962 436 974
rect 2 699 8 962
rect 38 954 48 962
rect 130 954 140 962
rect 174 960 310 962
rect 174 952 184 960
rect 80 934 90 944
rect 80 930 160 934
rect 208 930 218 942
rect 80 924 188 930
rect 130 916 140 924
rect 150 920 188 924
rect 208 920 264 930
rect 208 914 218 920
rect 38 900 48 906
rect 174 900 184 904
rect 14 890 184 900
rect 14 798 24 890
rect 300 872 310 960
rect 362 961 406 962
rect 362 954 367 961
rect 373 954 406 961
rect 362 952 406 954
rect 426 952 488 962
rect 426 946 436 952
rect 392 928 402 936
rect 337 927 402 928
rect 337 921 338 927
rect 344 921 402 927
rect 337 920 402 921
rect 38 869 310 872
rect 388 894 426 906
rect 438 894 468 906
rect 388 869 395 894
rect 38 862 395 869
rect 438 862 468 874
rect 38 854 48 862
rect 130 834 140 844
rect 186 852 196 862
rect 80 824 196 834
rect 278 832 288 842
rect 450 850 460 862
rect 450 840 543 850
rect 228 831 308 832
rect 228 824 300 831
rect 307 824 308 831
rect 450 830 460 840
rect 80 816 90 824
rect 228 822 308 824
rect 228 814 238 822
rect 442 818 470 830
rect 38 798 48 806
rect 130 798 140 806
rect 186 798 196 804
rect 278 798 288 804
rect 14 796 348 798
rect 14 791 97 796
rect 104 791 338 796
rect 14 789 338 791
rect 344 789 348 796
rect 14 788 348 789
rect 388 796 430 798
rect 388 790 394 796
rect 402 790 430 796
rect 388 786 430 790
rect 442 786 470 798
rect 741 721 807 731
rect 381 699 735 701
rect 2 691 735 699
rect 2 689 391 691
rect 119 681 129 689
rect 211 681 221 689
rect 305 675 315 689
rect 161 661 171 671
rect 161 653 241 661
rect 339 653 349 665
rect 161 651 319 653
rect 211 643 221 651
rect 231 643 319 651
rect 339 643 357 653
rect 339 637 349 643
rect 119 627 129 633
rect 95 624 241 627
rect 95 618 97 624
rect 104 621 241 624
rect 305 621 315 627
rect 104 618 315 621
rect 95 617 315 618
rect 95 606 105 617
rect 231 611 315 617
rect 95 600 96 606
rect 103 600 105 606
rect 95 473 105 600
rect 381 545 391 689
rect 463 683 473 691
rect 555 683 565 691
rect 649 677 659 691
rect 505 663 515 673
rect 505 655 585 663
rect 683 655 693 667
rect 505 653 663 655
rect 555 645 565 653
rect 575 645 663 653
rect 683 645 701 655
rect 683 639 693 645
rect 463 629 473 635
rect 119 535 391 545
rect 119 527 129 535
rect 211 527 221 535
rect 255 533 391 535
rect 255 525 265 533
rect 161 507 171 517
rect 161 503 241 507
rect 289 503 299 515
rect 161 497 269 503
rect 211 489 221 497
rect 231 493 269 497
rect 289 493 345 503
rect 289 487 299 493
rect 119 473 129 479
rect 255 473 265 477
rect 95 463 265 473
rect 95 371 105 463
rect 381 445 391 533
rect 119 435 391 445
rect 439 623 585 629
rect 649 623 659 629
rect 439 619 659 623
rect 439 475 449 619
rect 575 613 659 619
rect 725 625 735 691
rect 799 625 983 627
rect 797 617 983 625
rect 797 615 809 617
rect 725 547 735 615
rect 799 607 809 615
rect 973 613 983 617
rect 891 587 901 597
rect 1007 591 1017 603
rect 1029 591 1039 649
rect 911 587 987 591
rect 841 581 987 587
rect 1007 581 1039 591
rect 841 577 921 581
rect 841 569 851 577
rect 1007 575 1017 581
rect 463 537 735 547
rect 463 529 473 537
rect 555 529 565 537
rect 599 535 735 537
rect 599 527 609 535
rect 505 509 515 519
rect 505 505 585 509
rect 633 505 643 517
rect 505 499 613 505
rect 555 491 565 499
rect 575 495 613 499
rect 633 495 689 505
rect 633 489 643 495
rect 463 475 473 481
rect 599 475 609 479
rect 439 465 609 475
rect 119 427 129 435
rect 211 407 221 417
rect 267 425 277 435
rect 161 397 277 407
rect 359 405 369 415
rect 161 389 171 397
rect 309 395 379 405
rect 309 387 319 395
rect 119 371 129 379
rect 211 371 221 379
rect 267 371 277 377
rect 359 371 369 377
rect 439 373 449 465
rect 725 447 735 535
rect 463 437 735 447
rect 799 553 809 559
rect 891 553 901 559
rect 973 553 983 565
rect 799 543 983 553
rect 463 429 473 437
rect 555 409 565 419
rect 611 427 621 437
rect 505 399 621 409
rect 703 407 713 417
rect 505 391 515 399
rect 653 397 723 407
rect 653 389 663 397
rect 463 373 473 381
rect 555 373 565 381
rect 611 373 621 379
rect 703 373 713 379
rect 799 373 809 543
rect 921 541 983 543
rect 859 527 877 537
rect 439 371 809 373
rect 95 363 809 371
rect 95 361 449 363
<< metal2 >>
rect 151 1008 373 1013
rect 367 961 373 1008
rect 338 796 344 921
rect 97 624 104 791
rect 373 721 731 731
rect 373 653 383 721
rect 367 643 383 653
rect 701 537 711 645
rect 735 615 787 625
rect 701 527 849 537
rect 877 527 887 537
<< ntransistor >>
rect 412 936 416 946
rect 54 906 58 916
rect 122 906 126 916
rect 194 904 198 914
rect 426 882 438 886
rect 54 806 58 816
rect 122 806 126 816
rect 202 804 206 814
rect 270 804 274 814
rect 470 806 482 810
rect 135 633 139 643
rect 203 633 207 643
rect 325 627 329 637
rect 479 635 483 645
rect 547 635 551 645
rect 669 629 673 639
rect 815 559 819 569
rect 883 559 887 569
rect 993 565 997 575
rect 135 479 139 489
rect 203 479 207 489
rect 275 477 279 487
rect 479 481 483 491
rect 547 481 551 491
rect 619 479 623 489
rect 135 379 139 389
rect 203 379 207 389
rect 283 377 287 387
rect 351 377 355 387
rect 479 381 483 391
rect 547 381 551 391
rect 627 379 631 389
rect 695 379 699 389
<< ptransistor >>
rect 54 940 58 960
rect 122 940 126 960
rect 412 968 416 988
rect 194 936 198 956
rect 54 840 58 860
rect 122 840 126 860
rect 464 882 484 886
rect 202 838 206 858
rect 270 838 274 858
rect 426 806 446 810
rect 135 667 139 687
rect 203 667 207 687
rect 325 659 329 679
rect 479 669 483 689
rect 547 669 551 689
rect 669 661 673 681
rect 135 513 139 533
rect 203 513 207 533
rect 815 593 819 613
rect 883 593 887 613
rect 993 597 997 617
rect 275 509 279 529
rect 479 515 483 535
rect 547 515 551 535
rect 135 413 139 433
rect 203 413 207 433
rect 619 511 623 531
rect 283 411 287 431
rect 351 411 355 431
rect 479 415 483 435
rect 547 415 551 435
rect 627 413 631 433
rect 695 413 699 433
<< polycontact >>
rect 122 1008 127 1013
rect 12 965 19 970
rect 406 952 416 962
rect 488 952 498 962
rect 188 920 198 930
rect 264 920 274 930
rect 196 824 206 834
rect 300 824 307 831
rect 543 840 551 850
rect 394 790 402 796
rect 807 721 819 731
rect 319 643 329 653
rect 663 645 673 655
rect 96 600 103 606
rect 1029 649 1039 659
rect 987 581 997 591
rect 269 493 279 503
rect 345 493 355 503
rect 877 527 887 537
rect 613 495 623 505
rect 689 495 699 505
rect 277 397 287 407
rect 379 395 389 405
rect 621 399 631 409
rect 723 397 733 407
<< ndcontact >>
rect 392 936 402 946
rect 426 936 436 946
rect 38 906 48 916
rect 130 906 140 916
rect 174 904 184 914
rect 208 904 218 914
rect 426 894 438 906
rect 38 806 48 816
rect 80 806 90 816
rect 130 806 140 816
rect 186 804 196 814
rect 228 804 238 814
rect 278 804 288 814
rect 426 862 438 874
rect 470 818 482 830
rect 470 786 482 798
rect 119 633 129 643
rect 211 633 221 643
rect 305 627 315 637
rect 339 627 349 637
rect 463 635 473 645
rect 555 635 565 645
rect 649 629 659 639
rect 683 629 693 639
rect 799 559 809 569
rect 841 559 851 569
rect 891 559 901 569
rect 973 565 983 575
rect 1007 565 1017 575
rect 119 479 129 489
rect 211 479 221 489
rect 255 477 265 487
rect 289 477 299 487
rect 463 481 473 491
rect 555 481 565 491
rect 599 479 609 489
rect 633 479 643 489
rect 119 379 129 389
rect 161 379 171 389
rect 211 379 221 389
rect 267 377 277 387
rect 309 377 319 387
rect 359 377 369 387
rect 463 381 473 391
rect 505 381 515 391
rect 555 381 565 391
rect 611 379 621 389
rect 653 379 663 389
rect 703 379 713 389
<< pdcontact >>
rect 38 944 48 954
rect 80 944 90 954
rect 392 974 402 984
rect 426 974 436 984
rect 130 944 140 954
rect 174 942 184 952
rect 208 942 218 952
rect 38 844 48 854
rect 468 894 480 906
rect 130 844 140 854
rect 186 842 196 852
rect 278 842 288 852
rect 468 862 480 874
rect 430 818 442 830
rect 430 786 442 798
rect 119 671 129 681
rect 161 671 171 681
rect 211 671 221 681
rect 305 665 315 675
rect 339 665 349 675
rect 463 673 473 683
rect 505 673 515 683
rect 555 673 565 683
rect 649 667 659 677
rect 683 667 693 677
rect 119 517 129 527
rect 161 517 171 527
rect 799 597 809 607
rect 891 597 901 607
rect 973 603 983 613
rect 1007 603 1017 613
rect 211 517 221 527
rect 255 515 265 525
rect 289 515 299 525
rect 463 519 473 529
rect 505 519 515 529
rect 555 519 565 529
rect 599 517 609 527
rect 119 417 129 427
rect 633 517 643 527
rect 211 417 221 427
rect 267 415 277 425
rect 359 415 369 425
rect 463 419 473 429
rect 555 419 565 429
rect 611 417 621 427
rect 703 417 713 427
<< m2contact >>
rect 146 1008 151 1013
rect 367 954 373 961
rect 338 921 344 927
rect 97 791 104 796
rect 338 789 344 796
rect 731 721 741 731
rect 357 643 367 653
rect 97 618 104 624
rect 701 645 711 655
rect 725 615 735 625
rect 787 615 797 625
rect 849 527 859 537
<< labels >>
rlabel metal1 114 693 114 693 1 Vdd
rlabel polysilicon 1036 681 1036 681 7 Cout
rlabel polysilicon 136 745 136 745 5 Input1
rlabel polysilicon 745 403 745 403 1 Sum
rlabel metal1 300 792 300 792 1 GND
rlabel polycontact 302 826 302 826 1 Output
rlabel polysilicon 56 975 56 975 5 Input2
rlabel metal1 396 994 396 994 5 Vdd
rlabel metal1 396 922 396 922 1 GND
rlabel metal1 402 956 402 956 1 Ctrl
rlabel polysilicon 124 1015 124 1015 5 AbS
rlabel metal1 397 898 397 898 1 panw
rlabel polysilicon 549 797 549 797 1 MuxOut
rlabel polysilicon 397 780 397 780 1 Cin
rlabel polysilicon 16 975 16 975 1 Vdd
rlabel polysilicon 90 603 90 603 1 GND
<< end >>

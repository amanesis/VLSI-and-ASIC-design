magic
tech scmos
timestamp 1540495306
<< polysilicon >>
rect -46 44 -42 64
rect 22 44 26 64
rect -46 0 -42 24
rect 22 0 26 24
rect -46 -30 -42 -10
rect 22 -30 26 -10
<< ndiffusion >>
rect -64 -10 -62 0
rect -52 -10 -46 0
rect -42 -10 22 0
rect 26 -10 30 0
rect 40 -10 42 0
<< pdiffusion >>
rect -64 38 -46 44
rect -64 28 -62 38
rect -52 28 -46 38
rect -64 24 -46 28
rect -42 38 22 44
rect -42 28 -20 38
rect -10 28 22 38
rect -42 24 22 28
rect 26 38 42 44
rect 26 28 30 38
rect 40 28 42 38
rect 26 24 42 28
<< metal1 >>
rect -74 46 40 56
rect -62 38 -52 46
rect 30 38 40 46
rect -20 18 -10 28
rect -20 8 60 18
rect 30 0 40 8
rect -62 -16 -52 -10
rect -62 -26 60 -16
<< ntransistor >>
rect -46 -10 -42 0
rect 22 -10 26 0
<< ptransistor >>
rect -46 24 -42 44
rect 22 24 26 44
<< ndcontact >>
rect -62 -10 -52 0
rect 30 -10 40 0
<< pdcontact >>
rect -62 28 -52 38
rect -20 28 -10 38
rect 30 28 40 38
<< labels >>
rlabel metal1 54 12 54 12 1 Output
rlabel metal1 -72 50 -72 50 3 Vdd
rlabel metal1 52 -22 52 -22 1 GND
rlabel polysilicon -44 62 -44 62 5 Input1
rlabel polysilicon 24 61 24 61 5 Input2
<< end >>

magic
tech scmos
timestamp 1540545044
<< polysilicon >>
rect -270 166 -266 228
rect -202 166 -198 228
rect 74 168 78 188
rect 142 168 146 228
rect 410 210 414 212
rect 412 200 414 210
rect -80 158 -76 164
rect -270 122 -266 146
rect -202 122 -198 146
rect 264 160 268 166
rect -80 132 -76 138
rect 74 124 78 148
rect 142 124 146 148
rect 264 134 268 140
rect -80 116 -76 122
rect -270 12 -266 112
rect -202 12 -198 112
rect 264 118 268 124
rect -80 100 -76 106
rect -130 8 -126 28
rect 74 14 78 114
rect 142 14 146 114
rect 264 102 268 108
rect 410 92 414 200
rect 628 138 632 164
rect 478 92 482 112
rect 588 96 592 102
rect 410 48 414 72
rect 478 48 482 72
rect 588 70 592 76
rect 588 54 592 60
rect 588 38 592 44
rect -270 -32 -266 -8
rect -202 -32 -198 -8
rect 214 10 218 30
rect 410 18 414 38
rect 478 16 482 38
rect -130 -18 -126 -12
rect -54 -18 -50 -6
rect -130 -34 -126 -28
rect -270 -88 -266 -42
rect -202 -88 -198 -42
rect -130 -50 -126 -44
rect -122 -90 -118 -70
rect -54 -90 -50 -28
rect 74 -30 78 -6
rect 142 -30 146 -6
rect 478 4 482 6
rect 214 -16 218 -10
rect 290 -16 294 -4
rect 214 -32 218 -26
rect 74 -86 78 -40
rect 142 -86 146 -40
rect 214 -48 218 -42
rect -270 -132 -266 -108
rect -202 -132 -198 -108
rect 222 -88 226 -68
rect 290 -88 294 -26
rect -122 -114 -118 -110
rect -122 -134 -118 -124
rect -54 -134 -50 -110
rect 74 -118 78 -106
rect -16 -122 78 -118
rect 74 -130 78 -122
rect 142 -130 146 -106
rect 222 -112 226 -108
rect -270 -162 -266 -142
rect -202 -162 -198 -142
rect 222 -132 226 -122
rect 290 -132 294 -108
rect 328 -120 342 -116
rect -122 -164 -118 -144
rect -54 -164 -50 -144
rect 74 -160 78 -140
rect 142 -160 146 -140
rect 222 -162 226 -142
rect 290 -162 294 -142
<< ndiffusion >>
rect -288 112 -286 122
rect -276 112 -270 122
rect -266 112 -202 122
rect -198 112 -194 122
rect -184 112 -182 122
rect -102 106 -100 116
rect -90 106 -80 116
rect -76 106 -66 116
rect -56 106 -54 116
rect 56 114 58 124
rect 68 114 74 124
rect 78 114 142 124
rect 146 114 150 124
rect 160 114 162 124
rect 242 108 244 118
rect 254 108 264 118
rect 268 108 278 118
rect 288 108 290 118
rect 392 38 394 48
rect 404 38 410 48
rect 414 38 436 48
rect 446 38 478 48
rect 482 38 486 48
rect 496 38 498 48
rect 566 44 568 54
rect 578 44 588 54
rect 592 44 602 54
rect 612 44 614 54
rect -288 -42 -286 -32
rect -276 -42 -270 -32
rect -266 -42 -202 -32
rect -198 -42 -194 -32
rect -184 -42 -182 -32
rect -152 -44 -150 -34
rect -140 -44 -130 -34
rect -126 -44 -116 -34
rect -106 -44 -104 -34
rect 56 -40 58 -30
rect 68 -40 74 -30
rect 78 -40 142 -30
rect 146 -40 150 -30
rect 160 -40 162 -30
rect 192 -42 194 -32
rect 204 -42 214 -32
rect 218 -42 228 -32
rect 238 -42 240 -32
rect -288 -142 -286 -132
rect -276 -142 -270 -132
rect -266 -142 -244 -132
rect -234 -142 -202 -132
rect -198 -142 -194 -132
rect -184 -142 -182 -132
rect -140 -144 -138 -134
rect -128 -144 -122 -134
rect -118 -144 -96 -134
rect -86 -144 -54 -134
rect -50 -144 -46 -134
rect -36 -144 -34 -134
rect 56 -140 58 -130
rect 68 -140 74 -130
rect 78 -140 100 -130
rect 110 -140 142 -130
rect 146 -140 150 -130
rect 160 -140 162 -130
rect 204 -142 206 -132
rect 216 -142 222 -132
rect 226 -142 248 -132
rect 258 -142 290 -132
rect 294 -142 298 -132
rect 308 -142 310 -132
<< pdiffusion >>
rect -288 160 -270 166
rect -288 150 -286 160
rect -276 150 -270 160
rect -288 146 -270 150
rect -266 160 -202 166
rect -266 150 -244 160
rect -234 150 -202 160
rect -266 146 -202 150
rect -198 160 -182 166
rect -198 150 -194 160
rect -184 150 -182 160
rect 56 162 74 168
rect -198 146 -182 150
rect -102 154 -80 158
rect -102 144 -100 154
rect -90 144 -80 154
rect -102 138 -80 144
rect -76 154 -54 158
rect -76 144 -66 154
rect -56 144 -54 154
rect 56 152 58 162
rect 68 152 74 162
rect 56 148 74 152
rect 78 162 142 168
rect 78 152 100 162
rect 110 152 142 162
rect 78 148 142 152
rect 146 162 162 168
rect 146 152 150 162
rect 160 152 162 162
rect 146 148 162 152
rect 242 156 264 160
rect -76 138 -54 144
rect 242 146 244 156
rect 254 146 264 156
rect 242 140 264 146
rect 268 156 290 160
rect 268 146 278 156
rect 288 146 290 156
rect 268 140 290 146
rect -288 6 -270 12
rect -288 -4 -286 6
rect -276 -4 -270 6
rect -288 -8 -270 -4
rect -266 6 -202 12
rect -266 -4 -244 6
rect -234 -4 -202 6
rect -266 -8 -202 -4
rect -198 6 -182 12
rect 566 92 588 96
rect 392 86 410 92
rect 392 76 394 86
rect 404 76 410 86
rect 392 72 410 76
rect 414 72 478 92
rect 482 86 498 92
rect 482 76 486 86
rect 496 76 498 86
rect 566 82 568 92
rect 578 82 588 92
rect 566 76 588 82
rect 592 92 614 96
rect 592 82 602 92
rect 612 82 614 92
rect 592 76 614 82
rect 482 72 498 76
rect 56 8 74 14
rect -198 -4 -194 6
rect -184 -4 -182 6
rect -198 -8 -182 -4
rect -152 4 -130 8
rect -152 -6 -150 4
rect -140 -6 -130 4
rect -152 -12 -130 -6
rect -126 4 -104 8
rect -126 -6 -116 4
rect -106 -6 -104 4
rect 56 -2 58 8
rect 68 -2 74 8
rect 56 -6 74 -2
rect 78 8 142 14
rect 78 -2 100 8
rect 110 -2 142 8
rect 78 -6 142 -2
rect 146 8 162 14
rect 146 -2 150 8
rect 160 -2 162 8
rect 146 -6 162 -2
rect 192 6 214 10
rect 192 -4 194 6
rect 204 -4 214 6
rect -126 -12 -104 -6
rect -288 -94 -270 -88
rect -288 -104 -286 -94
rect -276 -104 -270 -94
rect -288 -108 -270 -104
rect -266 -108 -202 -88
rect -198 -94 -182 -88
rect 192 -10 214 -4
rect 218 6 240 10
rect 218 -4 228 6
rect 238 -4 240 6
rect 218 -10 240 -4
rect -198 -104 -194 -94
rect -184 -104 -182 -94
rect -198 -108 -182 -104
rect -140 -96 -122 -90
rect -140 -106 -138 -96
rect -128 -106 -122 -96
rect -140 -110 -122 -106
rect -118 -110 -54 -90
rect -50 -96 -34 -90
rect -50 -106 -46 -96
rect -36 -106 -34 -96
rect 56 -92 74 -86
rect 56 -102 58 -92
rect 68 -102 74 -92
rect 56 -106 74 -102
rect 78 -106 142 -86
rect 146 -92 162 -86
rect 146 -102 150 -92
rect 160 -102 162 -92
rect 146 -106 162 -102
rect 204 -94 222 -88
rect 204 -104 206 -94
rect 216 -104 222 -94
rect -50 -110 -34 -106
rect 204 -108 222 -104
rect 226 -108 290 -88
rect 294 -94 310 -88
rect 294 -104 298 -94
rect 308 -104 310 -94
rect 294 -108 310 -104
<< metal1 >>
rect 336 200 402 210
rect -24 178 330 180
rect -298 170 330 178
rect -298 168 -14 170
rect -286 160 -276 168
rect -194 160 -184 168
rect -100 154 -90 168
rect -244 140 -234 150
rect -244 132 -164 140
rect -66 132 -56 144
rect -244 130 -86 132
rect -194 122 -184 130
rect -174 122 -86 130
rect -66 122 -48 132
rect -66 116 -56 122
rect -286 106 -276 112
rect -310 100 -164 106
rect -100 100 -90 106
rect -310 96 -90 100
rect -310 -48 -300 96
rect -174 90 -90 96
rect -24 24 -14 168
rect 58 162 68 170
rect 150 162 160 170
rect 244 156 254 170
rect 100 142 110 152
rect 100 134 180 142
rect 278 134 288 146
rect 100 132 258 134
rect 150 124 160 132
rect 170 124 258 132
rect 278 124 296 134
rect 278 118 288 124
rect 58 108 68 114
rect -286 14 -14 24
rect -286 6 -276 14
rect -194 6 -184 14
rect -150 12 -14 14
rect -150 4 -140 12
rect -244 -14 -234 -4
rect -244 -18 -164 -14
rect -116 -18 -106 -6
rect -244 -24 -136 -18
rect -194 -32 -184 -24
rect -174 -28 -136 -24
rect -116 -28 -60 -18
rect -116 -34 -106 -28
rect -286 -48 -276 -42
rect -150 -48 -140 -44
rect -310 -58 -140 -48
rect -310 -150 -300 -58
rect -24 -76 -14 12
rect -286 -86 -14 -76
rect 34 102 180 108
rect 244 102 254 108
rect 34 98 254 102
rect 34 -46 44 98
rect 170 92 254 98
rect 320 104 330 170
rect 394 104 578 106
rect 392 96 578 104
rect 392 94 404 96
rect 320 26 330 94
rect 394 86 404 94
rect 568 92 578 96
rect 486 66 496 76
rect 602 70 612 82
rect 624 70 634 128
rect 506 66 582 70
rect 436 60 582 66
rect 602 60 634 70
rect 436 56 516 60
rect 436 48 446 56
rect 602 54 612 60
rect 58 16 330 26
rect 58 8 68 16
rect 150 8 160 16
rect 194 14 330 16
rect 194 6 204 14
rect 100 -12 110 -2
rect 100 -16 180 -12
rect 228 -16 238 -4
rect 100 -22 208 -16
rect 150 -30 160 -22
rect 170 -26 208 -22
rect 228 -26 284 -16
rect 228 -32 238 -26
rect 58 -46 68 -40
rect 194 -46 204 -42
rect 34 -56 204 -46
rect -286 -94 -276 -86
rect -194 -114 -184 -104
rect -138 -96 -128 -86
rect -244 -124 -128 -114
rect -46 -116 -36 -106
rect -244 -132 -234 -124
rect -96 -126 -26 -116
rect -96 -134 -86 -126
rect -286 -150 -276 -142
rect -194 -150 -184 -142
rect -138 -150 -128 -144
rect -46 -150 -36 -144
rect 34 -148 44 -56
rect 320 -74 330 14
rect 58 -84 330 -74
rect 394 32 404 38
rect 486 32 496 38
rect 568 32 578 44
rect 394 22 578 32
rect 58 -92 68 -84
rect 150 -112 160 -102
rect 206 -94 216 -84
rect 100 -122 216 -112
rect 298 -114 308 -104
rect 100 -130 110 -122
rect 248 -124 318 -114
rect 248 -132 258 -124
rect 58 -148 68 -140
rect 150 -148 160 -140
rect 206 -148 216 -142
rect 298 -148 308 -142
rect 394 -148 404 22
rect 516 20 578 22
rect 454 6 472 16
rect 34 -150 404 -148
rect -310 -158 404 -150
rect -310 -160 44 -158
<< metal2 >>
rect -32 200 326 210
rect -32 132 -22 200
rect -38 122 -22 132
rect 296 16 306 124
rect 330 94 382 104
rect 296 6 444 16
rect 472 6 482 16
<< ntransistor >>
rect -270 112 -266 122
rect -202 112 -198 122
rect -80 106 -76 116
rect 74 114 78 124
rect 142 114 146 124
rect 264 108 268 118
rect 410 38 414 48
rect 478 38 482 48
rect 588 44 592 54
rect -270 -42 -266 -32
rect -202 -42 -198 -32
rect -130 -44 -126 -34
rect 74 -40 78 -30
rect 142 -40 146 -30
rect 214 -42 218 -32
rect -270 -142 -266 -132
rect -202 -142 -198 -132
rect -122 -144 -118 -134
rect -54 -144 -50 -134
rect 74 -140 78 -130
rect 142 -140 146 -130
rect 222 -142 226 -132
rect 290 -142 294 -132
<< ptransistor >>
rect -270 146 -266 166
rect -202 146 -198 166
rect -80 138 -76 158
rect 74 148 78 168
rect 142 148 146 168
rect 264 140 268 160
rect -270 -8 -266 12
rect -202 -8 -198 12
rect 410 72 414 92
rect 478 72 482 92
rect 588 76 592 96
rect -130 -12 -126 8
rect 74 -6 78 14
rect 142 -6 146 14
rect -270 -108 -266 -88
rect -202 -108 -198 -88
rect 214 -10 218 10
rect -122 -110 -118 -90
rect -54 -110 -50 -90
rect 74 -106 78 -86
rect 142 -106 146 -86
rect 222 -108 226 -88
rect 290 -108 294 -88
<< polycontact >>
rect 402 200 412 210
rect -86 122 -76 132
rect 258 124 268 134
rect 624 128 634 138
rect 582 60 592 70
rect -136 -28 -126 -18
rect -60 -28 -50 -18
rect 472 6 482 16
rect 208 -26 218 -16
rect 284 -26 294 -16
rect -128 -124 -118 -114
rect -26 -126 -16 -116
rect 216 -122 226 -112
rect 318 -124 328 -114
<< ndcontact >>
rect -286 112 -276 122
rect -194 112 -184 122
rect -100 106 -90 116
rect -66 106 -56 116
rect 58 114 68 124
rect 150 114 160 124
rect 244 108 254 118
rect 278 108 288 118
rect 394 38 404 48
rect 436 38 446 48
rect 486 38 496 48
rect 568 44 578 54
rect 602 44 612 54
rect -286 -42 -276 -32
rect -194 -42 -184 -32
rect -150 -44 -140 -34
rect -116 -44 -106 -34
rect 58 -40 68 -30
rect 150 -40 160 -30
rect 194 -42 204 -32
rect 228 -42 238 -32
rect -286 -142 -276 -132
rect -244 -142 -234 -132
rect -194 -142 -184 -132
rect -138 -144 -128 -134
rect -96 -144 -86 -134
rect -46 -144 -36 -134
rect 58 -140 68 -130
rect 100 -140 110 -130
rect 150 -140 160 -130
rect 206 -142 216 -132
rect 248 -142 258 -132
rect 298 -142 308 -132
<< pdcontact >>
rect -286 150 -276 160
rect -244 150 -234 160
rect -194 150 -184 160
rect -100 144 -90 154
rect -66 144 -56 154
rect 58 152 68 162
rect 100 152 110 162
rect 150 152 160 162
rect 244 146 254 156
rect 278 146 288 156
rect -286 -4 -276 6
rect -244 -4 -234 6
rect 394 76 404 86
rect 486 76 496 86
rect 568 82 578 92
rect 602 82 612 92
rect -194 -4 -184 6
rect -150 -6 -140 4
rect -116 -6 -106 4
rect 58 -2 68 8
rect 100 -2 110 8
rect 150 -2 160 8
rect 194 -4 204 6
rect -286 -104 -276 -94
rect 228 -4 238 6
rect -194 -104 -184 -94
rect -138 -106 -128 -96
rect -46 -106 -36 -96
rect 58 -102 68 -92
rect 150 -102 160 -92
rect 206 -104 216 -94
rect 298 -104 308 -94
<< m2contact >>
rect 326 200 336 210
rect -48 122 -38 132
rect 296 124 306 134
rect 320 94 330 104
rect 382 94 392 104
rect 444 6 454 16
<< labels >>
rlabel metal1 -291 172 -291 172 1 Vdd
rlabel metal1 -304 100 -304 100 1 GND
rlabel polysilicon 144 225 144 225 5 Cin
rlabel polysilicon 631 160 631 160 7 Cout
rlabel polysilicon -269 224 -269 224 5 Input1
rlabel polysilicon -200 224 -200 224 5 Input2
rlabel polysilicon 340 -118 340 -118 1 Sum
<< end >>

magic
tech scmos
timestamp 1540495531
<< polysilicon >>
rect 28 74 32 94
rect 96 74 100 94
rect 28 30 32 54
rect 96 30 100 54
rect 28 0 32 20
rect 96 0 100 20
<< ndiffusion >>
rect 10 20 12 30
rect 22 20 28 30
rect 32 20 54 30
rect 64 20 96 30
rect 100 20 104 30
rect 114 20 116 30
<< pdiffusion >>
rect 10 68 28 74
rect 10 58 12 68
rect 22 58 28 68
rect 10 54 28 58
rect 32 54 96 74
rect 100 68 116 74
rect 100 58 104 68
rect 114 58 116 68
rect 100 54 116 58
<< metal1 >>
rect 0 76 22 86
rect 12 68 22 76
rect 104 48 114 58
rect 54 38 134 48
rect 54 30 64 38
rect 12 14 22 20
rect 104 14 114 20
rect 12 4 134 14
<< ntransistor >>
rect 28 20 32 30
rect 96 20 100 30
<< ptransistor >>
rect 28 54 32 74
rect 96 54 100 74
<< ndcontact >>
rect 12 20 22 30
rect 54 20 64 30
rect 104 20 114 30
<< pdcontact >>
rect 12 58 22 68
rect 104 58 114 68
<< labels >>
rlabel metal1 128 42 128 42 1 Output
rlabel metal1 2 80 2 80 3 Vdd
rlabel metal1 126 8 126 8 1 GND
rlabel polysilicon 30 93 30 93 5 Input1
rlabel polysilicon 98 92 98 92 5 Input2
<< end >>

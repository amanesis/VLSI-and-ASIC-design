magic
tech scmos
timestamp 1542285287
<< polysilicon >>
rect 6 30 16 32
rect 6 6 16 10
rect 6 -14 16 -10
rect 6 -26 16 -24
<< ndiffusion >>
rect -20 -24 -18 -14
rect -8 -24 6 -14
rect 16 -24 28 -14
rect 38 -24 40 -14
<< pdiffusion >>
rect -20 26 6 30
rect -20 16 -18 26
rect -8 16 6 26
rect -20 10 6 16
rect 16 26 40 30
rect 16 16 28 26
rect 38 16 40 26
rect 16 10 40 16
<< metal1 >>
rect 6 42 16 50
rect -18 4 -8 16
rect -26 -6 -8 4
rect -18 -14 -8 -6
rect 28 4 38 16
rect 28 -6 46 4
rect 28 -14 38 -6
<< ntransistor >>
rect 6 -24 16 -14
<< ptransistor >>
rect 6 10 16 30
<< polycontact >>
rect 6 32 16 42
rect 6 -36 16 -26
<< ndcontact >>
rect -18 -24 -8 -14
rect 28 -24 38 -14
<< pdcontact >>
rect -18 16 -8 26
rect 28 16 38 26
<< labels >>
rlabel metal1 -24 0 -24 0 3 Input
rlabel metal1 42 0 42 0 7 Output
rlabel metal1 10 46 10 46 5 C
<< end >>

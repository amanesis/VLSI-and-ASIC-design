magic
tech scmos
timestamp 1543680363
<< polysilicon >>
rect 7736 680 7747 683
rect 68 651 72 655
rect 68 546 72 646
rect 408 630 414 633
rect 250 606 254 609
rect 4551 574 4561 587
rect 1506 483 1516 520
rect 3028 506 3038 534
rect 4320 436 4325 457
rect -39 339 -33 344
rect 25 314 33 320
rect 1558 310 1563 314
rect 3081 310 3086 314
rect 20 205 33 212
rect 4578 175 4586 673
rect 7736 673 7738 680
rect 7745 673 7747 680
rect 6299 651 6303 654
rect 6077 551 6087 583
rect 6299 546 6303 646
rect 7736 554 7747 673
rect 7737 483 7747 554
rect 9259 506 9269 576
rect 10782 574 10792 614
rect 12308 568 12323 575
rect 12308 551 12318 568
rect 6077 424 6087 427
rect 6077 418 6079 424
rect 6085 418 6087 424
rect 6077 416 6087 418
rect 6194 339 6201 344
rect 4603 311 4612 320
rect 6259 314 6264 320
rect 7789 310 7794 314
rect 9312 309 9317 314
rect 10834 310 10843 320
rect 6238 206 6239 212
rect 6246 206 6264 212
rect 6238 205 6264 206
rect 4578 168 4603 175
rect 10824 168 10834 175
rect 626 -20 630 -10
<< metal1 >>
rect 4586 673 7738 680
rect 73 646 6298 651
rect 4985 625 6640 630
rect 4825 601 6481 606
rect 6085 418 6141 424
rect 6201 344 6208 346
rect 6201 206 6208 339
rect 6239 212 6246 223
rect 6035 196 6059 206
rect 6070 196 6208 206
rect 5729 -10 6857 -4
<< metal2 >>
rect 6008 476 6332 482
rect 6008 426 6015 476
rect 6326 424 6332 476
rect 6141 229 6147 418
rect 6141 223 6239 229
<< polycontact >>
rect 4578 673 4586 680
rect 68 646 73 651
rect 7738 673 7745 680
rect 6298 646 6303 651
rect 6079 418 6085 424
rect 6201 339 6208 344
rect 6239 206 6246 212
<< m2contact >>
rect 6008 420 6015 426
rect 6141 418 6147 424
rect 6326 418 6332 424
rect 6239 223 6246 229
use Register_4Bit  Register_4Bit_0
timestamp 1543589226
transform 1 0 103 0 1 67
box -136 -77 5984 563
use Register_4Bit  Register_4Bit_1
timestamp 1543589226
transform 1 0 6334 0 1 67
box -136 -77 5984 563
<< labels >>
rlabel polysilicon 7742 550 7742 550 1 Out3
rlabel polysilicon 9264 575 9264 575 1 Out2
rlabel polysilicon 10787 610 10787 610 1 Out1
rlabel polysilicon 4556 583 4556 583 1 Out5
rlabel polysilicon 3033 529 3033 529 1 Out6
rlabel polysilicon 1511 514 1511 514 1 Out7
rlabel polysilicon 4323 453 4323 453 1 Vdd
rlabel polysilicon 25 208 25 208 1 SR
rlabel polysilicon 10829 171 10829 171 1 SL
rlabel polysilicon 628 -16 628 -16 1 CLK
rlabel polysilicon 10838 312 10838 312 1 In0
rlabel polysilicon 9314 312 9314 312 1 In1
rlabel polysilicon 7791 312 7791 312 1 In2
rlabel polysilicon 6261 317 6261 317 1 In3
rlabel polysilicon 4607 313 4607 313 1 In4
rlabel polysilicon 3083 312 3083 312 1 In5
rlabel polysilicon 1560 312 1560 312 1 In6
rlabel polysilicon 27 317 27 317 1 In7
rlabel polysilicon 6081 578 6081 578 1 Out4
rlabel polysilicon 411 632 411 632 5 CLR
rlabel polysilicon 252 608 252 608 1 Ctrl1
rlabel polysilicon 70 653 70 653 1 Ctrl0
rlabel polysilicon 12320 571 12320 571 7 Out0
rlabel polysilicon 6196 342 6196 342 1 GND
<< end >>

magic
tech scmos
timestamp 1543586722
<< polysilicon >>
rect 504 425 510 435
rect 330 405 336 413
rect 1197 392 1202 395
rect -10 364 -6 370
rect 172 365 176 371
rect -10 338 -6 344
rect 72 338 76 354
rect 172 339 176 345
rect 254 339 258 355
rect -30 330 -25 336
rect 1428 339 1438 349
rect -10 322 -6 328
rect -42 273 -34 279
rect -10 262 -6 312
rect 72 262 76 328
rect 172 323 176 329
rect -10 258 4 262
rect 16 258 20 262
rect 38 258 42 262
rect 62 258 76 262
rect -10 186 -6 258
rect 72 186 76 258
rect -10 182 4 186
rect 24 182 28 186
rect 44 182 48 186
rect 60 182 76 186
rect 172 263 176 313
rect 254 263 258 329
rect 505 322 509 331
rect 1428 319 1438 329
rect 505 307 509 314
rect 172 259 186 263
rect 198 259 202 263
rect 220 259 224 263
rect 244 259 258 263
rect 172 187 176 259
rect 254 187 258 259
rect 172 183 186 187
rect 206 183 210 187
rect 226 183 230 187
rect 242 183 258 187
rect -42 164 -34 171
rect -40 127 -34 134
rect -10 115 -6 182
rect 72 115 76 182
rect 548 134 552 193
rect 646 156 650 187
rect 646 134 650 140
rect 1076 134 1080 187
rect 548 126 552 129
rect 646 126 650 129
rect 1076 125 1080 129
rect -10 111 4 115
rect 16 111 21 115
rect 36 111 42 115
rect 62 111 76 115
rect -10 29 -6 111
rect 72 29 76 111
rect -10 25 4 29
rect 24 25 28 29
rect 46 25 50 29
rect 62 25 76 29
rect -43 9 -37 15
<< ndiffusion >>
rect -32 312 -30 322
rect -20 312 -10 322
rect -6 312 4 322
rect 14 312 16 322
rect 4 282 16 284
rect 4 262 16 270
rect 150 313 152 323
rect 162 313 172 323
rect 176 313 186 323
rect 196 313 198 323
rect 4 250 16 258
rect 4 236 16 238
rect 48 206 60 208
rect 48 186 60 194
rect 186 283 198 285
rect 186 263 198 271
rect 186 251 198 259
rect 186 237 198 239
rect 230 207 242 209
rect 230 187 242 195
rect 48 174 60 182
rect 48 160 60 162
rect 4 136 16 138
rect 4 115 16 124
rect 230 175 242 183
rect 230 161 242 163
rect 4 104 16 111
rect 4 90 16 92
rect 50 50 62 52
rect 50 29 62 38
rect 50 18 62 25
rect 50 4 62 6
<< pdiffusion >>
rect -32 360 -10 364
rect -32 350 -30 360
rect -20 350 -10 360
rect -32 344 -10 350
rect -6 360 16 364
rect -6 350 4 360
rect 14 350 16 360
rect 150 361 172 365
rect -6 344 16 350
rect 150 351 152 361
rect 162 351 172 361
rect 150 345 172 351
rect 176 361 198 365
rect 176 351 186 361
rect 196 351 198 361
rect 176 345 198 351
rect 42 282 62 284
rect 42 270 46 282
rect 58 270 62 282
rect 42 262 62 270
rect 42 250 62 258
rect 42 238 46 250
rect 58 238 62 250
rect 42 236 62 238
rect 4 206 24 208
rect 4 194 8 206
rect 20 194 24 206
rect 4 186 24 194
rect 224 283 244 285
rect 224 271 228 283
rect 240 271 244 283
rect 224 263 244 271
rect 224 251 244 259
rect 224 239 228 251
rect 240 239 244 251
rect 224 237 244 239
rect 186 207 206 209
rect 186 195 190 207
rect 202 195 206 207
rect 186 187 206 195
rect 4 174 24 182
rect 4 162 8 174
rect 20 162 24 174
rect 4 160 24 162
rect 42 136 62 138
rect 42 124 46 136
rect 58 124 62 136
rect 42 115 62 124
rect 186 175 206 183
rect 186 163 190 175
rect 202 163 206 175
rect 186 161 206 163
rect 42 104 62 111
rect 42 92 46 104
rect 58 92 62 104
rect 42 90 62 92
rect 4 50 24 52
rect 4 38 8 50
rect 20 38 24 50
rect 4 29 24 38
rect 4 18 24 25
rect 4 6 8 18
rect 20 6 24 18
rect 4 4 24 6
<< metal1 >>
rect 152 417 418 425
rect 152 384 162 417
rect 310 409 322 417
rect 520 411 644 421
rect 520 409 574 411
rect 634 387 644 411
rect 764 387 774 389
rect 1194 387 1197 389
rect 1202 387 1204 389
rect -30 375 162 384
rect -30 360 -20 375
rect 152 361 162 375
rect 302 363 319 373
rect 366 369 430 379
rect 626 377 700 387
rect 710 377 1130 387
rect 1140 377 1368 387
rect 364 363 370 369
rect 536 363 572 373
rect 608 363 610 375
rect 4 338 14 350
rect 186 339 196 351
rect -22 336 -16 338
rect -19 330 -16 336
rect -22 328 -16 330
rect 4 328 66 338
rect 160 329 166 339
rect 186 329 248 339
rect 312 329 430 339
rect 542 335 566 345
rect 4 322 14 328
rect 186 323 196 329
rect -30 304 -20 312
rect 152 304 162 313
rect -30 296 277 304
rect -34 279 4 282
rect -28 273 4 279
rect -34 270 4 273
rect 16 270 46 282
rect 138 271 186 283
rect 198 271 228 283
rect 16 238 46 250
rect 28 226 38 238
rect 138 226 148 271
rect 198 239 228 251
rect 28 216 148 226
rect 210 227 220 239
rect 294 227 302 315
rect 210 217 302 227
rect 468 304 482 335
rect 498 314 503 322
rect 468 296 471 304
rect 478 296 482 304
rect 28 206 38 216
rect 210 207 220 217
rect 20 194 48 206
rect 202 195 230 207
rect 468 177 482 296
rect 626 271 636 377
rect 840 375 850 377
rect 928 375 938 377
rect 528 261 636 271
rect 626 255 636 261
rect 682 361 774 371
rect 584 219 594 225
rect 682 219 692 361
rect 804 329 848 339
rect 896 329 936 339
rect 984 329 998 339
rect 764 269 774 285
rect 764 219 774 259
rect 584 209 634 219
rect 692 209 708 219
rect 756 209 774 219
rect 804 213 814 329
rect 840 287 928 297
rect 980 213 990 329
rect 1056 255 1066 377
rect 1270 375 1280 377
rect 1358 375 1368 377
rect 1112 361 1204 371
rect 804 203 826 213
rect 898 203 990 213
rect 1112 219 1122 361
rect 1234 329 1278 339
rect 1326 329 1366 339
rect 1414 329 1428 339
rect 1194 269 1204 285
rect 1194 219 1204 259
rect 1122 209 1138 219
rect 1186 209 1204 219
rect 1234 213 1244 329
rect 1270 287 1358 297
rect 1410 213 1420 329
rect 1234 203 1256 213
rect 1328 203 1420 213
rect 1410 197 1420 203
rect 528 177 538 183
rect -34 171 8 174
rect -28 164 8 171
rect -34 162 8 164
rect 20 162 48 174
rect 142 163 190 175
rect 202 163 230 175
rect 468 167 710 177
rect 700 165 710 167
rect -34 134 4 136
rect -27 127 4 134
rect -34 125 4 127
rect 16 124 46 136
rect 16 92 46 104
rect 28 75 37 92
rect 142 75 154 163
rect 700 155 826 165
rect 858 149 868 173
rect 946 167 1140 177
rect 946 165 956 167
rect 888 155 928 165
rect 938 155 956 165
rect 1130 165 1140 167
rect 1130 155 1256 165
rect 1288 149 1298 173
rect 1318 155 1358 165
rect 1368 155 1386 165
rect 1410 155 1421 165
rect 553 129 645 134
rect 650 129 1075 134
rect 28 67 154 75
rect 28 50 37 67
rect 20 38 50 50
rect -37 15 8 18
rect -31 9 8 15
rect -37 6 8 9
rect 20 6 50 18
rect -25 -15 -15 6
rect 1410 -15 1420 135
rect -25 -22 1420 -15
<< metal2 >>
rect 668 395 732 409
rect 668 375 680 395
rect 620 363 680 375
rect 302 315 492 322
rect 294 314 492 315
rect 285 296 471 304
rect 700 265 710 377
rect 722 325 732 395
rect 998 403 1162 413
rect 998 339 1008 403
rect 774 259 858 269
rect 682 149 692 209
rect 928 165 938 287
rect 1130 265 1140 377
rect 1152 325 1162 403
rect 1204 259 1288 269
rect 836 155 878 165
rect 1112 149 1122 209
rect 1358 165 1368 287
rect 1266 155 1308 165
rect 682 139 858 149
rect 1112 139 1288 149
rect 1410 145 1420 186
<< ntransistor >>
rect -10 312 -6 322
rect 172 313 176 323
rect 4 258 16 262
rect 48 182 60 186
rect 186 259 198 263
rect 230 183 242 187
rect 4 111 16 115
rect 50 25 62 29
<< ptransistor >>
rect -10 344 -6 364
rect 172 345 176 365
rect 42 258 62 262
rect 4 182 24 186
rect 224 259 244 263
rect 186 183 206 187
rect 42 111 62 115
rect 4 25 24 29
<< polycontact >>
rect 1197 387 1202 392
rect 430 369 442 379
rect -25 330 -19 336
rect -16 328 -6 338
rect 66 328 76 338
rect 166 329 176 339
rect 248 329 258 339
rect -34 273 -28 279
rect 503 314 509 322
rect 1428 329 1438 339
rect -34 164 -28 171
rect -34 127 -27 134
rect 548 129 553 134
rect 645 129 650 134
rect 1075 129 1080 134
rect -37 9 -31 15
<< ndcontact >>
rect -30 312 -20 322
rect 4 312 14 322
rect 4 270 16 282
rect 152 313 162 323
rect 186 313 196 323
rect 4 238 16 250
rect 48 194 60 206
rect 186 271 198 283
rect 186 239 198 251
rect 230 195 242 207
rect 48 162 60 174
rect 4 124 16 136
rect 230 163 242 175
rect 4 92 16 104
rect 50 38 62 50
rect 50 6 62 18
<< pdcontact >>
rect -30 350 -20 360
rect 4 350 14 360
rect 152 351 162 361
rect 186 351 196 361
rect 46 270 58 282
rect 46 238 58 250
rect 8 194 20 206
rect 228 271 240 283
rect 228 239 240 251
rect 190 195 202 207
rect 8 162 20 174
rect 46 124 58 136
rect 190 163 202 175
rect 46 92 58 104
rect 8 38 20 50
rect 8 6 20 18
<< m2contact >>
rect 700 377 710 387
rect 1130 377 1140 387
rect 610 363 620 375
rect 294 315 302 322
rect 277 296 285 304
rect 492 314 498 322
rect 471 296 478 304
rect 998 329 1008 339
rect 722 315 732 325
rect 700 255 710 265
rect 764 259 774 269
rect 682 209 692 219
rect 928 287 938 297
rect 858 259 868 269
rect 1152 315 1162 325
rect 1130 255 1140 265
rect 1194 259 1204 269
rect 1112 209 1122 219
rect 1358 287 1368 297
rect 1288 259 1298 269
rect 1410 186 1420 197
rect 826 155 836 165
rect 878 155 888 165
rect 928 155 938 165
rect 1256 155 1266 165
rect 858 139 868 149
rect 1308 155 1318 165
rect 1358 155 1368 165
rect 1288 139 1298 149
rect 1410 135 1420 145
use Inverter  Inverter_10
timestamp 1540453251
transform 1 0 347 0 1 339
box -38 -8 20 70
use NAND  NAND_0
timestamp 1540495306
transform 1 0 483 0 1 361
box -74 -30 60 64
use Inverter  Inverter_9
timestamp 1540453251
transform 1 0 600 0 1 340
box -38 -8 20 70
use gate  gate_0
timestamp 1542285287
transform 1 0 758 0 1 321
box -26 -36 46 50
use Inverter  Inverter_2
timestamp 1540453251
transform 1 0 876 0 1 305
box -38 -8 20 70
use Inverter  Inverter_3
timestamp 1540453251
transform 1 0 964 0 1 305
box -38 -8 20 70
use gate  gate_2
timestamp 1542285287
transform 1 0 1188 0 1 321
box -26 -36 46 50
use Inverter  Inverter_4
timestamp 1540453251
transform 1 0 1306 0 1 305
box -38 -8 20 70
use Inverter  Inverter_5
timestamp 1540453251
transform 1 0 1394 0 1 305
box -38 -8 20 70
use Inverter  Inverter_8
timestamp 1540453251
transform 1 0 564 0 1 191
box -38 -8 20 70
use Inverter  Inverter_0
timestamp 1540453251
transform 1 0 662 0 1 185
box -38 -8 20 70
use Inverter  Inverter_1
timestamp 1540453251
transform 1 0 736 0 1 185
box -38 -8 20 70
use gate  gate_1
timestamp 1542285287
transform 1 0 852 0 1 209
box -26 -36 46 50
use Inverter  Inverter_6
timestamp 1540453251
transform 1 0 1092 0 1 185
box -38 -8 20 70
use Inverter  Inverter_7
timestamp 1540453251
transform 1 0 1166 0 1 185
box -38 -8 20 70
use gate  gate_3
timestamp 1542285287
transform 1 0 1282 0 1 209
box -26 -36 46 50
<< labels >>
rlabel metal1 -26 298 -26 298 1 GND
rlabel metal1 156 299 156 299 1 GND
rlabel metal1 950 159 950 159 1 GND
rlabel polysilicon 1434 345 1434 345 7 Q
rlabel metal1 1380 159 1380 159 1 GND
rlabel polysilicon 508 431 508 431 5 D
rlabel polysilicon 332 409 332 409 1 CLR
rlabel metal1 163 334 163 334 1 ctrl1
rlabel polysilicon -28 333 -28 333 1 Ctrl0
rlabel polysilicon -39 277 -39 277 3 Input1
rlabel polysilicon -39 167 -39 167 3 Input2
rlabel polysilicon -37 130 -37 130 3 Input3
rlabel polysilicon -40 12 -40 12 3 Input4
rlabel polysilicon 1200 394 1200 394 1 Vdd
rlabel polysilicon 550 127 550 127 1 CLK
<< end >>

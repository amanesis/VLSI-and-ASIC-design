magic
tech scmos
timestamp 1543589226
<< polysilicon >>
rect 305 558 306 563
rect -35 344 -31 474
rect 147 345 151 534
rect 305 387 311 558
rect 1827 558 1828 563
rect 1449 505 1452 506
rect 1449 497 1451 505
rect 1172 369 1177 413
rect 1403 323 1413 416
rect -136 272 -54 277
rect -70 247 -67 253
rect 502 191 509 196
rect -70 138 -67 145
rect -59 108 -52 114
rect 523 -71 527 153
rect 621 -71 625 84
rect 1051 -71 1055 127
rect 1449 108 1452 497
rect 1487 454 1491 474
rect 1487 344 1491 449
rect 1669 345 1673 534
rect 1827 387 1833 558
rect 3350 558 3351 563
rect 2969 484 2975 487
rect 2969 477 2972 484
rect 2925 437 2935 439
rect 2925 323 2935 428
rect 1455 253 1460 256
rect 1449 101 1459 108
rect 2045 -71 2049 153
rect 2143 -71 2147 83
rect 2573 -71 2577 127
rect 2969 108 2975 477
rect 3010 344 3014 449
rect 3192 345 3196 534
rect 3350 387 3356 558
rect 4876 558 4877 563
rect 4448 505 4458 507
rect 4456 497 4458 505
rect 4448 323 4458 497
rect 4536 344 4540 449
rect 4718 345 4722 534
rect 4876 387 4882 558
rect 5974 478 5976 484
rect 5982 478 5984 484
rect 5974 323 5984 478
rect 2978 253 2983 256
rect 4500 253 4509 256
rect 2969 101 2980 108
rect 3568 -71 3572 153
rect 3666 -71 3670 87
rect 4096 -71 4100 127
rect 4500 101 4506 108
rect 5094 -71 5098 153
rect 5192 -71 5196 88
rect 5622 -71 5626 127
<< metal1 >>
rect 311 558 1828 563
rect 1833 558 3351 563
rect 3356 558 4877 563
rect 152 534 1668 539
rect 1673 534 3191 539
rect 3196 534 4717 539
rect 1459 497 4448 505
rect -31 474 1486 479
rect 2979 478 5976 484
rect 5982 478 5984 484
rect 2979 477 5984 478
rect 1492 449 3009 454
rect 3014 449 4535 454
rect -119 428 2925 437
rect -119 110 -110 428
rect 1343 351 1473 361
rect 2865 351 2995 361
rect 4388 351 4526 361
rect 1424 270 1467 278
rect 2950 270 2990 278
rect 4476 270 4516 278
rect -53 139 -50 145
rect 1424 139 1434 270
rect 1463 148 1470 150
rect 2950 139 2958 270
rect 2991 247 2998 254
rect 2986 148 2994 150
rect 4476 139 4488 270
rect 4516 248 4523 254
rect 4512 148 4520 150
rect 1361 129 1385 139
rect 1395 129 1434 139
rect 2883 129 2958 139
rect 4406 128 4488 139
rect -119 99 -59 110
rect 4515 101 4523 108
rect 529 -77 619 -71
rect 627 -77 1049 -71
rect 1058 -77 2043 -71
rect 2049 -77 2140 -71
rect 2150 -77 2570 -71
rect 2580 -77 3566 -71
rect 3572 -77 3662 -71
rect 3673 -77 4092 -71
rect 4104 -77 5092 -71
rect 5098 -77 5189 -71
rect 5200 -77 5619 -71
<< metal2 >>
rect 1385 150 1463 157
rect 2907 152 2986 157
rect 2917 150 2986 152
rect 4430 150 4512 157
<< polycontact >>
rect 306 558 311 563
rect 147 534 152 539
rect -35 474 -31 479
rect 1828 558 1833 563
rect 1668 534 1673 539
rect 1451 497 1459 505
rect -54 272 -49 277
rect 509 191 514 196
rect 1486 474 1491 479
rect 1487 449 1492 454
rect 3351 558 3356 563
rect 3191 534 3196 539
rect 2972 477 2979 484
rect 2925 428 2935 437
rect 3009 449 3014 454
rect 4877 558 4882 563
rect 4717 534 4722 539
rect 4448 497 4456 505
rect 4535 449 4540 454
rect 5976 478 5982 484
rect 523 -77 529 -71
rect 619 -77 627 -71
rect 1049 -77 1058 -71
rect 2043 -77 2049 -71
rect 2140 -77 2150 -71
rect 2570 -77 2580 -71
rect 3566 -77 3572 -71
rect 3662 -77 3673 -71
rect 4092 -77 4104 -71
rect 5092 -77 5098 -71
rect 5189 -77 5200 -71
rect 5619 -77 5626 -71
<< m2contact >>
rect 1385 160 1395 171
rect 1463 150 1470 157
rect 2986 150 2994 157
rect 4512 150 4520 157
use Mux_D_Flip_Fop  Mux_D_Flip_Fop_0
timestamp 1543586722
transform 1 0 -25 0 1 -26
box -43 -22 1438 435
use Mux_D_Flip_Fop  Mux_D_Flip_Fop_1
timestamp 1543586722
transform 1 0 1497 0 1 -26
box -43 -22 1438 435
use Mux_D_Flip_Fop  Mux_D_Flip_Fop_2
timestamp 1543586722
transform 1 0 3020 0 1 -26
box -43 -22 1438 435
use Mux_D_Flip_Fop  Mux_D_Flip_Fop_3
timestamp 1543586722
transform 1 0 4546 0 1 -26
box -43 -22 1438 435
<< labels >>
rlabel space 285 292 285 292 1 MuxOut
rlabel space 619 343 619 343 1 NandOut
rlabel space 781 294 781 294 1 LatchOut
rlabel space 969 308 969 308 1 QOut
rlabel polysilicon -68 142 -68 142 1 SR
rlabel polysilicon -69 250 -69 250 1 In3
rlabel polysilicon 1457 254 1457 254 1 In2
rlabel polysilicon 2980 255 2980 255 1 In1
rlabel polysilicon -33 471 -33 471 1 Ctrl0
rlabel polysilicon 308 544 308 544 1 CLR
rlabel polysilicon 149 504 149 504 1 Ctrl1
rlabel polysilicon 4501 255 4501 255 1 In0
rlabel polysilicon 4501 105 4501 105 1 SL
rlabel polysilicon 4452 424 4452 424 1 Out1
rlabel polysilicon 5979 428 5979 428 7 Out0
rlabel polysilicon 2930 421 2930 421 1 Out2
rlabel polysilicon 1408 413 1408 413 1 Out3
rlabel polysilicon 525 -61 525 -61 1 CLK
rlabel polysilicon 1174 412 1174 412 1 Vdd
rlabel polysilicon -128 274 -128 274 1 GND
<< end >>

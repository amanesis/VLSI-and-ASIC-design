magic
tech scmos
timestamp 1540498033
<< polysilicon >>
rect 8 278 12 298
rect 76 278 80 298
rect 198 270 202 276
rect 8 234 12 258
rect 76 234 80 258
rect 198 244 202 250
rect 198 228 202 234
rect 8 124 12 224
rect 76 124 80 224
rect 198 212 202 218
rect 148 120 152 140
rect 8 80 12 104
rect 76 80 80 104
rect 148 94 152 100
rect 224 94 228 106
rect 148 78 152 84
rect 8 24 12 70
rect 76 24 80 70
rect 148 62 152 68
rect 156 22 160 42
rect 224 22 228 84
rect 8 -20 12 4
rect 76 -20 80 4
rect 156 -2 160 2
rect 156 -22 160 -12
rect 224 -22 228 2
rect 262 -10 310 -6
rect 8 -50 12 -30
rect 76 -50 80 -30
rect 156 -52 160 -32
rect 224 -52 228 -32
<< ndiffusion >>
rect -10 224 -8 234
rect 2 224 8 234
rect 12 224 76 234
rect 80 224 84 234
rect 94 224 96 234
rect 176 218 178 228
rect 188 218 198 228
rect 202 218 212 228
rect 222 218 224 228
rect -10 70 -8 80
rect 2 70 8 80
rect 12 70 76 80
rect 80 70 84 80
rect 94 70 96 80
rect 126 68 128 78
rect 138 68 148 78
rect 152 68 162 78
rect 172 68 174 78
rect -10 -30 -8 -20
rect 2 -30 8 -20
rect 12 -30 34 -20
rect 44 -30 76 -20
rect 80 -30 84 -20
rect 94 -30 96 -20
rect 138 -32 140 -22
rect 150 -32 156 -22
rect 160 -32 182 -22
rect 192 -32 224 -22
rect 228 -32 232 -22
rect 242 -32 244 -22
<< pdiffusion >>
rect -10 272 8 278
rect -10 262 -8 272
rect 2 262 8 272
rect -10 258 8 262
rect 12 272 76 278
rect 12 262 34 272
rect 44 262 76 272
rect 12 258 76 262
rect 80 272 96 278
rect 80 262 84 272
rect 94 262 96 272
rect 80 258 96 262
rect 176 266 198 270
rect 176 256 178 266
rect 188 256 198 266
rect 176 250 198 256
rect 202 266 224 270
rect 202 256 212 266
rect 222 256 224 266
rect 202 250 224 256
rect -10 118 8 124
rect -10 108 -8 118
rect 2 108 8 118
rect -10 104 8 108
rect 12 118 76 124
rect 12 108 34 118
rect 44 108 76 118
rect 12 104 76 108
rect 80 118 96 124
rect 80 108 84 118
rect 94 108 96 118
rect 80 104 96 108
rect 126 116 148 120
rect 126 106 128 116
rect 138 106 148 116
rect 126 100 148 106
rect 152 116 174 120
rect 152 106 162 116
rect 172 106 174 116
rect 152 100 174 106
rect -10 18 8 24
rect -10 8 -8 18
rect 2 8 8 18
rect -10 4 8 8
rect 12 4 76 24
rect 80 18 96 24
rect 80 8 84 18
rect 94 8 96 18
rect 80 4 96 8
rect 138 16 156 22
rect 138 6 140 16
rect 150 6 156 16
rect 138 2 156 6
rect 160 2 224 22
rect 228 16 244 22
rect 228 6 232 16
rect 242 6 244 16
rect 228 2 244 6
<< metal1 >>
rect -20 280 264 290
rect -8 272 2 280
rect 84 272 94 280
rect 178 266 188 280
rect 34 252 44 262
rect 34 244 114 252
rect 212 244 222 256
rect 34 242 192 244
rect 84 234 94 242
rect 104 234 192 242
rect 212 234 234 244
rect 212 228 222 234
rect -8 218 2 224
rect -32 212 114 218
rect 178 212 188 218
rect -32 208 188 212
rect -32 64 -22 208
rect 104 202 188 208
rect 254 136 264 280
rect -8 126 264 136
rect -8 118 2 126
rect 84 118 94 126
rect 128 124 264 126
rect 128 116 138 124
rect 34 98 44 108
rect 34 94 114 98
rect 162 94 172 106
rect 34 88 142 94
rect 84 80 94 88
rect 104 84 142 88
rect 162 84 218 94
rect 162 78 172 84
rect -8 64 2 70
rect 128 64 138 68
rect -32 54 138 64
rect -32 -38 -22 54
rect 254 36 264 124
rect -8 26 264 36
rect -8 18 2 26
rect 84 -2 94 8
rect 140 16 150 26
rect 34 -12 150 -2
rect 232 -4 242 6
rect 34 -20 44 -12
rect 182 -14 250 -4
rect 182 -22 192 -14
rect -8 -38 2 -30
rect 84 -38 94 -30
rect 140 -38 150 -32
rect 232 -38 242 -32
rect -32 -48 262 -38
<< ntransistor >>
rect 8 224 12 234
rect 76 224 80 234
rect 198 218 202 228
rect 8 70 12 80
rect 76 70 80 80
rect 148 68 152 78
rect 8 -30 12 -20
rect 76 -30 80 -20
rect 156 -32 160 -22
rect 224 -32 228 -22
<< ptransistor >>
rect 8 258 12 278
rect 76 258 80 278
rect 198 250 202 270
rect 8 104 12 124
rect 76 104 80 124
rect 148 100 152 120
rect 8 4 12 24
rect 76 4 80 24
rect 156 2 160 22
rect 224 2 228 22
<< polycontact >>
rect 192 234 202 244
rect 142 84 152 94
rect 218 84 228 94
rect 150 -12 160 -2
rect 250 -14 262 -4
<< ndcontact >>
rect -8 224 2 234
rect 84 224 94 234
rect 178 218 188 228
rect 212 218 222 228
rect -8 70 2 80
rect 84 70 94 80
rect 128 68 138 78
rect 162 68 172 78
rect -8 -30 2 -20
rect 34 -30 44 -20
rect 84 -30 94 -20
rect 140 -32 150 -22
rect 182 -32 192 -22
rect 232 -32 242 -22
<< pdcontact >>
rect -8 262 2 272
rect 34 262 44 272
rect 84 262 94 272
rect 178 256 188 266
rect 212 256 222 266
rect -8 108 2 118
rect 34 108 44 118
rect 84 108 94 118
rect 128 106 138 116
rect 162 106 172 116
rect -8 8 2 18
rect 84 8 94 18
rect 140 6 150 16
rect 232 6 242 16
<< labels >>
rlabel metal1 -15 285 -15 285 1 Vdd
rlabel polysilicon 10 296 10 296 5 Input1
rlabel polysilicon 78 295 78 295 5 Input2
rlabel metal1 253 -45 253 -45 1 GND
rlabel metal1 228 238 228 238 1 Cout
rlabel polysilicon 301 -8 301 -8 1 Sum
<< end >>
